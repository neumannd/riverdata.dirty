netcdf river40_1 {
dimensions:
	longitude = 1 ;
	latitude = 1 ;
	depth = 1 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float longitude(longitude) ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:axis = "X" ;
	float latitude(latitude) ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:axis = "Y" ;
	float depth(depth) ;
		depth:units = "m" ;
		depth:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:units = "day as %Y%m%d.%f" ;
		time:calendar = "proleptic_gregorian" ;
	float mole_concentration_of_ammonium_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_ammonium_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_ammonium_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_ammonium_in_seawater:standard_name = "mole_concentration_of_ammonium_in_seawater";
	float mole_concentration_of_nitrate_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_nitrate_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_nitrate_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_nitrate_in_seawater:standard_name = "mole_concentration_of_nitrate_in_seawater" ;
	float mole_concentration_of_phosphate_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_phosphate_in_seawater:units = "mmol P/m3" ;
		mole_concentration_of_phosphate_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_phosphate_in_seawater:standard_name = "mole_concentration_of_phosphate_in_seawater" ;
	float mole_concentration_of_diatoms_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_diatoms_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_diatoms_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_diatoms_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_diatoms_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_flagellates_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_flagellates_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_flagellates_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_flagellates_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_flagellates_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_cyanobacteria_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_cyanobacteria_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_cyanobacteria_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_cyanobacteria_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_cyanobacteria_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_zooplankton_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_zooplankton_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_zooplankton_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_zooplankton_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_zooplankton_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_detritus_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_detritus_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_detritus_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_detritus_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_detritus_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_oxygen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_oxygen_in_seawater:units = "mmol O/m3" ;
		mole_concentration_of_oxygen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_oxygen_in_seawater:standard_name = "mole_concentration_of_oxygen_in_seawater" ;
	float mole_concentration_of_silicate_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_silicate_in_seawater:units = "mmol Si/m3" ;
		mole_concentration_of_silicate_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_silicate_in_seawater:standard_name = "mole_concentration_of_silicate_in_seawater" ;
	float mole_concentration_of_protozooplankton_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_protozooplankton_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_protozooplankton_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_protozooplankton_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_protozooplankton_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_detritus_expressed_as_silicate_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_detritus_expressed_as_silicate_in_seawater:units = "mmol Si/m3" ;
		mole_concentration_of_detritus_expressed_as_silicate_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_detritus_expressed_as_silicate_in_seawater:standard_name = "mole_concentration_of_detritus_expressed_as_silicate_in_seawater" ;
	float mole_concentration_of_labile_dissolved_organic_nitrogen_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_labile_dissolved_organic_nitrogen_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_ammonium_from_warnow_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_ammonium_from_warnow_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_ammonium_from_warnow_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_ammonium_from_warnow_in_seawater:standard_name = "mole_concentration_of_ammonium_from_warnow_in_seawater";
	float mole_concentration_of_nitrate_from_warnow_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_nitrate_from_warnow_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_nitrate_from_warnow_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_nitrate_from_warnow_in_seawater:standard_name = "mole_concentration_of_nitrate_from_warnow_in_seawater" ;
	float mole_concentration_of_phosphate_from_warnow_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_phosphate_from_warnow_in_seawater:units = "mmol P/m3" ;
		mole_concentration_of_phosphate_from_warnow_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_phosphate_from_warnow_in_seawater:standard_name = "mole_concentration_of_phosphate_from_warnow_in_seawater" ;
	float mole_concentration_of_diatoms_from_warnow_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_diatoms_from_warnow_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_diatoms_from_warnow_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_diatoms_from_warnow_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_diatoms_from_warnow_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_flagellates_from_warnow_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_flagellates_from_warnow_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_flagellates_from_warnow_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_flagellates_from_warnow_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_flagellates_from_warnow_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_cyanobacteria_from_warnow_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_cyanobacteria_from_warnow_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_cyanobacteria_from_warnow_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_cyanobacteria_from_warnow_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_cyanobacteria_from_warnow_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_zooplankton_from_warnow_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_zooplankton_from_warnow_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_zooplankton_from_warnow_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_zooplankton_from_warnow_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_zooplankton_from_warnow_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_detritus_from_warnow_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_detritus_from_warnow_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_detritus_from_warnow_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_detritus_from_warnow_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_detritus_from_warnow_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_oxygen_from_warnow_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_oxygen_from_warnow_in_seawater:units = "mmol O/m3" ;
		mole_concentration_of_oxygen_from_warnow_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_oxygen_from_warnow_in_seawater:standard_name = "mole_concentration_of_oxygen_from_warnow_in_seawater" ;
	float mole_concentration_of_silicate_from_warnow_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_silicate_from_warnow_in_seawater:units = "mmol Si/m3" ;
		mole_concentration_of_silicate_from_warnow_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_silicate_from_warnow_in_seawater:standard_name = "mole_concentration_of_silicate_from_warnow_in_seawater" ;
	float mole_concentration_of_protozooplankton_from_warnow_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_protozooplankton_from_warnow_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_protozooplankton_from_warnow_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_protozooplankton_from_warnow_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_protozooplankton_from_warnow_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_detritus_from_warnow_expressed_as_silicate_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_detritus_from_warnow_expressed_as_silicate_in_seawater:units = "mmol Si/m3" ;
		mole_concentration_of_detritus_from_warnow_expressed_as_silicate_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_detritus_from_warnow_expressed_as_silicate_in_seawater:standard_name = "mole_concentration_of_detritus_from_warnow_expressed_as_silicate_in_seawater" ;
	float mole_concentration_of_labile_dissolved_organic_nitrogen_from_warnow_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_from_warnow_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_from_warnow_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_from_warnow_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_labile_dissolved_organic_nitrogen_from_warnow_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_ammonium_from_trave_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_ammonium_from_trave_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_ammonium_from_trave_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_ammonium_from_trave_in_seawater:standard_name = "mole_concentration_of_ammonium_from_trave_in_seawater";
	float mole_concentration_of_nitrate_from_trave_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_nitrate_from_trave_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_nitrate_from_trave_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_nitrate_from_trave_in_seawater:standard_name = "mole_concentration_of_nitrate_from_trave_in_seawater" ;
	float mole_concentration_of_phosphate_from_trave_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_phosphate_from_trave_in_seawater:units = "mmol P/m3" ;
		mole_concentration_of_phosphate_from_trave_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_phosphate_from_trave_in_seawater:standard_name = "mole_concentration_of_phosphate_from_trave_in_seawater" ;
	float mole_concentration_of_diatoms_from_trave_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_diatoms_from_trave_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_diatoms_from_trave_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_diatoms_from_trave_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_diatoms_from_trave_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_flagellates_from_trave_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_flagellates_from_trave_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_flagellates_from_trave_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_flagellates_from_trave_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_flagellates_from_trave_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_cyanobacteria_from_trave_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_cyanobacteria_from_trave_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_cyanobacteria_from_trave_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_cyanobacteria_from_trave_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_cyanobacteria_from_trave_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_zooplankton_from_trave_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_zooplankton_from_trave_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_zooplankton_from_trave_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_zooplankton_from_trave_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_zooplankton_from_trave_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_detritus_from_trave_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_detritus_from_trave_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_detritus_from_trave_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_detritus_from_trave_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_detritus_from_trave_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_oxygen_from_trave_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_oxygen_from_trave_in_seawater:units = "mmol O/m3" ;
		mole_concentration_of_oxygen_from_trave_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_oxygen_from_trave_in_seawater:standard_name = "mole_concentration_of_oxygen_from_trave_in_seawater" ;
	float mole_concentration_of_silicate_from_trave_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_silicate_from_trave_in_seawater:units = "mmol Si/m3" ;
		mole_concentration_of_silicate_from_trave_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_silicate_from_trave_in_seawater:standard_name = "mole_concentration_of_silicate_from_trave_in_seawater" ;
	float mole_concentration_of_protozooplankton_from_trave_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_protozooplankton_from_trave_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_protozooplankton_from_trave_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_protozooplankton_from_trave_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_protozooplankton_from_trave_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_detritus_from_trave_expressed_as_silicate_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_detritus_from_trave_expressed_as_silicate_in_seawater:units = "mmol Si/m3" ;
		mole_concentration_of_detritus_from_trave_expressed_as_silicate_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_detritus_from_trave_expressed_as_silicate_in_seawater:standard_name = "mole_concentration_of_detritus_from_trave_expressed_as_silicate_in_seawater" ;
	float mole_concentration_of_labile_dissolved_organic_nitrogen_from_trave_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_from_trave_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_from_trave_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_from_trave_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_labile_dissolved_organic_nitrogen_from_trave_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_ammonium_from_peene_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_ammonium_from_peene_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_ammonium_from_peene_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_ammonium_from_peene_in_seawater:standard_name = "mole_concentration_of_ammonium_from_peene_in_seawater";
	float mole_concentration_of_nitrate_from_peene_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_nitrate_from_peene_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_nitrate_from_peene_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_nitrate_from_peene_in_seawater:standard_name = "mole_concentration_of_nitrate_from_peene_in_seawater" ;
	float mole_concentration_of_phosphate_from_peene_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_phosphate_from_peene_in_seawater:units = "mmol P/m3" ;
		mole_concentration_of_phosphate_from_peene_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_phosphate_from_peene_in_seawater:standard_name = "mole_concentration_of_phosphate_from_peene_in_seawater" ;
	float mole_concentration_of_diatoms_from_peene_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_diatoms_from_peene_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_diatoms_from_peene_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_diatoms_from_peene_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_diatoms_from_peene_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_flagellates_from_peene_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_flagellates_from_peene_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_flagellates_from_peene_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_flagellates_from_peene_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_flagellates_from_peene_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_cyanobacteria_from_peene_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_cyanobacteria_from_peene_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_cyanobacteria_from_peene_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_cyanobacteria_from_peene_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_cyanobacteria_from_peene_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_zooplankton_from_peene_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_zooplankton_from_peene_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_zooplankton_from_peene_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_zooplankton_from_peene_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_zooplankton_from_peene_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_detritus_from_peene_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_detritus_from_peene_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_detritus_from_peene_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_detritus_from_peene_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_detritus_from_peene_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_oxygen_from_peene_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_oxygen_from_peene_in_seawater:units = "mmol O/m3" ;
		mole_concentration_of_oxygen_from_peene_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_oxygen_from_peene_in_seawater:standard_name = "mole_concentration_of_oxygen_from_peene_in_seawater" ;
	float mole_concentration_of_silicate_from_peene_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_silicate_from_peene_in_seawater:units = "mmol Si/m3" ;
		mole_concentration_of_silicate_from_peene_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_silicate_from_peene_in_seawater:standard_name = "mole_concentration_of_silicate_from_peene_in_seawater" ;
	float mole_concentration_of_protozooplankton_from_peene_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_protozooplankton_from_peene_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_protozooplankton_from_peene_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_protozooplankton_from_peene_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_protozooplankton_from_peene_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_detritus_from_peene_expressed_as_silicate_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_detritus_from_peene_expressed_as_silicate_in_seawater:units = "mmol Si/m3" ;
		mole_concentration_of_detritus_from_peene_expressed_as_silicate_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_detritus_from_peene_expressed_as_silicate_in_seawater:standard_name = "mole_concentration_of_detritus_from_peene_expressed_as_silicate_in_seawater" ;
	float mole_concentration_of_labile_dissolved_organic_nitrogen_from_peene_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_from_peene_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_from_peene_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_from_peene_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_labile_dissolved_organic_nitrogen_from_peene_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_ammonium_from_schwentine_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_ammonium_from_schwentine_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_ammonium_from_schwentine_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_ammonium_from_schwentine_in_seawater:standard_name = "mole_concentration_of_ammonium_from_schwentine_in_seawater";
	float mole_concentration_of_nitrate_from_schwentine_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_nitrate_from_schwentine_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_nitrate_from_schwentine_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_nitrate_from_schwentine_in_seawater:standard_name = "mole_concentration_of_nitrate_from_schwentine_in_seawater" ;
	float mole_concentration_of_phosphate_from_schwentine_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_phosphate_from_schwentine_in_seawater:units = "mmol P/m3" ;
		mole_concentration_of_phosphate_from_schwentine_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_phosphate_from_schwentine_in_seawater:standard_name = "mole_concentration_of_phosphate_from_schwentine_in_seawater" ;
	float mole_concentration_of_diatoms_from_schwentine_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_diatoms_from_schwentine_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_diatoms_from_schwentine_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_diatoms_from_schwentine_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_diatoms_from_schwentine_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_flagellates_from_schwentine_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_flagellates_from_schwentine_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_flagellates_from_schwentine_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_flagellates_from_schwentine_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_flagellates_from_schwentine_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_cyanobacteria_from_schwentine_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_cyanobacteria_from_schwentine_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_cyanobacteria_from_schwentine_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_cyanobacteria_from_schwentine_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_cyanobacteria_from_schwentine_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_zooplankton_from_schwentine_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_zooplankton_from_schwentine_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_zooplankton_from_schwentine_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_zooplankton_from_schwentine_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_zooplankton_from_schwentine_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_detritus_from_schwentine_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_detritus_from_schwentine_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_detritus_from_schwentine_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_detritus_from_schwentine_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_detritus_from_schwentine_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_oxygen_from_schwentine_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_oxygen_from_schwentine_in_seawater:units = "mmol O/m3" ;
		mole_concentration_of_oxygen_from_schwentine_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_oxygen_from_schwentine_in_seawater:standard_name = "mole_concentration_of_oxygen_from_schwentine_in_seawater" ;
	float mole_concentration_of_silicate_from_schwentine_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_silicate_from_schwentine_in_seawater:units = "mmol Si/m3" ;
		mole_concentration_of_silicate_from_schwentine_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_silicate_from_schwentine_in_seawater:standard_name = "mole_concentration_of_silicate_from_schwentine_in_seawater" ;
	float mole_concentration_of_protozooplankton_from_schwentine_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_protozooplankton_from_schwentine_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_protozooplankton_from_schwentine_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_protozooplankton_from_schwentine_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_protozooplankton_from_schwentine_expressed_as_nitrogen_in_seawater" ;
	float mole_concentration_of_detritus_from_schwentine_expressed_as_silicate_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_detritus_from_schwentine_expressed_as_silicate_in_seawater:units = "mmol Si/m3" ;
		mole_concentration_of_detritus_from_schwentine_expressed_as_silicate_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_detritus_from_schwentine_expressed_as_silicate_in_seawater:standard_name = "mole_concentration_of_detritus_from_schwentine_expressed_as_silicate_in_seawater" ;
	float mole_concentration_of_labile_dissolved_organic_nitrogen_from_schwentine_expressed_as_nitrogen_in_seawater(time, depth, latitude, longitude) ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_from_schwentine_expressed_as_nitrogen_in_seawater:units = "mmol N/m3" ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_from_schwentine_expressed_as_nitrogen_in_seawater:river_name = "RIVERNAME" ;
		mole_concentration_of_labile_dissolved_organic_nitrogen_from_schwentine_expressed_as_nitrogen_in_seawater:standard_name = "mole_concentration_of_labile_dissolved_organic_nitrogen_from_schwentine_expressed_as_nitrogen_in_seawater" ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:standard_name_vocabulary = "CF Standard Names 1.6";
		:history = "" ;
		:contact = "Thomas Neumann";
		:contact_email = "thomas.neumann@hzg.de";
		:originator = "Daniel Neumann";
		:contributor_name = "Thomas Neumann";
		:institution = "Leibniz Institute for Baltic Sea Research Warnemuende, Rostock-Warnemuende, Germany";
		:source = "compiled from MOM input";
		:summary = "River inflow into the southern Baltic Sea.";
		:title = "River inflow into the southern Baltic Sea.";
    :creationTime = "2017-06-19T12:00:00Z";
		:date_created = "2017-06-19";
		:date_modified = "2017-06-19";
    
data:

 mole_concentration_of_ammonium_in_seawater = 0.f, 0.f ;
 mole_concentration_of_nitrate_in_seawater = 0.f, 0.f ;
 mole_concentration_of_phosphate_in_seawater = 0.f, 0.f ;
 mole_concentration_of_diatoms_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_flagellates_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_cyanobacteria_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_zooplankton_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_detritus_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_oxygen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_silicate_in_seawater = 0.f, 0.f ;
 mole_concentration_of_protozooplankton_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_detritus_expressed_as_silicate_in_seawater = 0.f, 0.f ;
 mole_concentration_of_labile_dissolved_organic_nitrogen_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_ammonium_from_warnow_in_seawater = 0.f, 0.f ;
 mole_concentration_of_nitrate_from_warnow_in_seawater = 0.f, 0.f ;
 mole_concentration_of_phosphate_from_warnow_in_seawater = 0.f, 0.f ;
 mole_concentration_of_diatoms_from_warnow_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_flagellates_from_warnow_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_cyanobacteria_from_warnow_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_zooplankton_from_warnow_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_detritus_from_warnow_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_oxygen_from_warnow_in_seawater = 0.f, 0.f ;
 mole_concentration_of_silicate_from_warnow_in_seawater = 0.f, 0.f ;
 mole_concentration_of_protozooplankton_from_warnow_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_detritus_from_warnow_expressed_as_silicate_in_seawater = 0.f, 0.f ;
 mole_concentration_of_labile_dissolved_organic_nitrogen_from_warnow_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_ammonium_from_trave_in_seawater = 0.f, 0.f ;
 mole_concentration_of_nitrate_from_trave_in_seawater = 0.f, 0.f ;
 mole_concentration_of_phosphate_from_trave_in_seawater = 0.f, 0.f ;
 mole_concentration_of_diatoms_from_trave_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_flagellates_from_trave_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_cyanobacteria_from_trave_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_zooplankton_from_trave_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_detritus_from_trave_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_oxygen_from_trave_in_seawater = 0.f, 0.f ;
 mole_concentration_of_silicate_from_trave_in_seawater = 0.f, 0.f ;
 mole_concentration_of_protozooplankton_from_trave_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_detritus_from_trave_expressed_as_silicate_in_seawater = 0.f, 0.f ;
 mole_concentration_of_labile_dissolved_organic_nitrogen_from_trave_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_ammonium_from_peene_in_seawater = 0.f, 0.f ;
 mole_concentration_of_nitrate_from_peene_in_seawater = 0.f, 0.f ;
 mole_concentration_of_phosphate_from_peene_in_seawater = 0.f, 0.f ;
 mole_concentration_of_diatoms_from_peene_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_flagellates_from_peene_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_cyanobacteria_from_peene_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_zooplankton_from_peene_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_detritus_from_peene_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_oxygen_from_peene_in_seawater = 0.f, 0.f ;
 mole_concentration_of_silicate_from_peene_in_seawater = 0.f, 0.f ;
 mole_concentration_of_protozooplankton_from_peene_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_detritus_from_peene_expressed_as_silicate_in_seawater = 0.f, 0.f ;
 mole_concentration_of_labile_dissolved_organic_nitrogen_from_peene_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_ammonium_from_schwentine_in_seawater = 0.f, 0.f ;
 mole_concentration_of_nitrate_from_schwentine_in_seawater = 0.f, 0.f ;
 mole_concentration_of_phosphate_from_schwentine_in_seawater = 0.f, 0.f ;
 mole_concentration_of_diatoms_from_schwentine_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_flagellates_from_schwentine_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_cyanobacteria_from_schwentine_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_zooplankton_from_schwentine_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_detritus_from_schwentine_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_oxygen_from_schwentine_in_seawater = 0.f, 0.f ;
 mole_concentration_of_silicate_from_schwentine_in_seawater = 0.f, 0.f ;
 mole_concentration_of_protozooplankton_from_schwentine_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
 mole_concentration_of_detritus_from_schwentine_expressed_as_silicate_in_seawater = 0.f, 0.f ;
 mole_concentration_of_labile_dissolved_organic_nitrogen_from_schwentine_expressed_as_nitrogen_in_seawater = 0.f, 0.f ;
}